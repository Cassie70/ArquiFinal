library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity ROM_RGB is port(
	clk: in std_logic;
	clr: in std_logic;
	address: in std_logic_vector(7 downto 0);
	data_out : out std_logic_vector(23 downto 0)
);
end ROM_RGB;

architecture a_ROM_RGB of ROM_RGB is
	
	type ROM_Array is array (0 to 255) of std_logic_vector(23 downto 0);
	constant content: ROM_Array := (
		--1
		0=>"000000001110011111100111",
		1=>"010101001101010110000001",
		2=>"001010101010101110000001",
		3=>"010101000101010000000000",
		4=>"001010100010101000000000",
		5=>"010101001101010110000001",
		6=>"001010101010101110000001",
		7=>"000000001110011111100111",
		--2
		8=>"000000001111111111111111",
		9=>"000000001000000110000001",
		10=>"000000001000000110000001",
		11=>"000000000000000000000000",
		12=>"000000000000000000000000",
		13=>"000000001000000110000001",
		14=>"000000001000000110000001",
		15=>"000000001111111111111111",
		--3
		16=>"000000001111111111111111",
		17=>"000000001000000110000001",
		18=>"000000001011110110000001",
		19=>"000000001010010010000000",
		20=>"000000001010010010000000",
		21=>"000000001011110110000001",
		22=>"000000001000000110000001",
		23=>"000000001110011111100111",
		--4
		24=>"000000001110011111100111",
		25=>"000000001000000110000001",
		26=>"000000001000000110000001",
		27=>"000000001000000110000001",
		28=>"000000001000000110000001",
		29=>"000000001000000110000001",
		30=>"000000001000000110000001",
		31=>"000000001111111111111111",
		--5
		32=>"000000001111111111111111",
		33=>"000000001000000110010001",
		34=>"000000001000000110001101",
		35=>"000000000000000000111110",
		36=>"000000000000000000111110",
		37=>"000000001000000110001101",
		38=>"000000001000000110010001",
		39=>"000000001111111111111111",
		--6
		40=>"000000001111111111111111",
		41=>"011111101000000110000001",
		42=>"000000001000000110000001",
		43=>"000000000000000000000000",
		44=>"000000000000000000000000",
		45=>"000000001000000110000001",
		46=>"011111101000000110000001",
		47=>"000000001111111111111111",
		--7
		48=>"000000001110011111100111",
		49=>"000000001000000110000001",
		50=>"001001001000000110100101",
		51=>"001001000000000100100101",
		52=>"000000000000000100000001",
		53=>"000110001000000110011001",
		54=>"000000001000000110000001",
		55=>"000000001110011111100111",
		--8
		56=>"000000001111111111100111",
		57=>"000000001111111110000001",
		58=>"000000001111111110000001",
		59=>"000000001111111110000001",
		60=>"000000001111111110000001",
		61=>"000000001111111110000001",
		62=>"000000001111111110000001",
		63=>"000000001111111111100111",
		--9
		64=>"000110001110011111111111",
		65=>"011111101000000111111111",
		66=>"011111101000000111111111",
		67=>"111111100000000111111111",
		68=>"111111100000000111111111",
		69=>"011111101000000111111111",
		70=>"011111101000000111111111",
		71=>"000000001111111111111111",
		--10
		72=>"000110001110011111100111",
		73=>"011110001000000110000111",
		74=>"011111001000000110000011",
		75=>"011111101000000110000001",
		76=>"011101101000100110000001",
		77=>"011111101000000111111111",
		78=>"011111101110000110011111",
		79=>"000110001110011111111111",
		--11
		80=>"000000001111111111111111",
		81=>"011111101110011111111111",
		82=>"011111101110011111111111",
		83=>"111111110001100011111111",
		84=>"111111110011110011111111",
		85=>"011111101011110111111111",
		86=>"011111101010010111111111",
		87=>"000000001111111111111111",
		--12 animacion 1 FUEGOO
		88=>"111111111111111111111111",
		89=>"111111111111111111111111",
		90=>"110111101111111111111111",
		91=>"100010001101111011111111",
		92=>"100000001101110011111111",
		93=>"000000001000000011111110",
		94=>"000000000000000011001100",
		95=>"000000000000000010000100",
		--12 animacion 2
		96=>"111110111111111111111111",
		97=>"111110111111111111111111",
		98=>"001100011111101111111111",
		99=>"001000000111101111111111",
		100=>"000000000010000111111111",
		101=>"000000000000000001111011",
		102=>"000000000000000001111001",
		103=>"000000000000000001010000",
		--12 animacion 3
		104=>"111111111111111111111111",
		105=>"111111111111111111111111",
		106=>"111111011111111111111111",
		107=>"110110001111110111111111",
		108=>"100000001101110111111111",
		109=>"000000001001000011111111",
		110=>"000000000000000001111011",
		111=>"000000000000000000100001",
		--12 animacion 4
		112=>"111111111111111111111111",
		113=>"111111111111111111111111",
		114=>"111111111111111111111111",
		115=>"111011111111111111111111",
		116=>"110001101110111111111111",
		117=>"110000001110011011111111",
		118=>"000000001100010011101111",
		119=>"000000000000000011000110",
		--12 animacion 5
		120=>"111011111111111111111111",
		121=>"110001111110111111111111",
		122=>"100001111110111111111111",
		123=>"000000011000011111111111",
		124=>"000000001000000111101111",
		125=>"000000000000000011001111",
		126=>"000000000000000011000111",
		127=>"000000000000000010000010",
		--13 animacion 1 CARITA
		128=>"110000111100001111111111",
		129=>"100000011000000111111111",
		130=>"001001000010010011111111",
		131=>"001001000010010011111111",
		132=>"000000000000000011111111",
		133=>"010000100100001011111111",
		134=>"001111000011110011111111",
		135=>"100000011000000111111111",
		--14 animacion 2
		136=>"111111111100001111000011",
		137=>"111111111000000110000001",
		138=>"111111110010010000100100",
		139=>"111111110010010000100100",
		140=>"111111110000000000000000",
		141=>"111111110001100000011000",
		142=>"111111110010010000100100",
		143=>"111111111000000110000001",
		--14 animacion 3
		144=>"110000111111111111111111",
		145=>"100000011111111111111111",
		146=>"010000101111111111111111",
		147=>"001001001111111111111111",
		148=>"000000001111111111111111",
		149=>"000110001111111111111111",
		150=>"001111001111111111111111",
		151=>"100000011111111111111111",
		--15 animacion 1 corazon uwu
		152=>"000000001111111100000000",
		153=>"011001101111111101100110",
		154=>"100110011011111110111111",
		155=>"100000011011111110111111",
		156=>"100000011011111110111111",
		157=>"010000101101111101011110",
		158=>"001001001110011100100100",
		159=>"000110001111111100011000",
		--15 animacion 2
		160=>"000000000000000011111111",
		161=>"011001100110011011111111",
		162=>"100110011101111111011111",
		163=>"100000011100011111000111",
		164=>"100000011111001111110011",
		165=>"010000100111101011111011",
		166=>"001001000011110011111111",
		167=>"000110000001100011111111",
		--15 animacion 3
		168=>"111111110000000000000000",
		169=>"111111110110011001100110",
		170=>"100110011111100111111001",
		171=>"100000011111110111111101",
		172=>"100000011111111111111111",
		173=>"110000110111111001111110",
		174=>"111001110011110000111100",
		175=>"111111110001100000011000",
		--16 animacion 1 gei
		176=>"111111111111111111111111",
		177=>"111111111111111111111111",
		178=>"001111111111111111111111",
		179=>"001111110011111111111111",
		180=>"111111110011111111111111",
		181=>"111111111111111100111111",
		182=>"001111111111111100111111",
		183=>"111111111111111111111111",
		--16 animacion 2
		184=>"111111111111111111111111",
		185=>"111111111111111111111111",
		186=>"000011111111111111111111",
		187=>"000011110000111111111111",
		188=>"111111110000111111111111",
		189=>"111111111111111100001111",
		190=>"000011111111111100001111",
		191=>"111111111111111111111111",
		--16 animacion 3
		192=>"111111111111111111111111",
		193=>"111111111111111111111111",
		194=>"000000001111111111111111",
		195=>"000000000000000011111111",
		196=>"111111110000000011111111",
		197=>"111111111111111100000000",
		198=>"000000001111111100000000",
		199=>"111111111111111111111111",
		--16 animacion 4
		200=>"111111111111111111111111",
		201=>"111111111111111111111111",
		202=>"111111110000000000000000",
		203=>"000000001111111100000000",
		204=>"000000000000000000000000",
		205=>"000000001111111100000000",
		206=>"111111110000000000000000",
		207=>"111111111111111111111111",
		others => x"FFFFFF"
	);
begin
	process(clk,clr,address)
	begin
		if(clr='1') then	
			data_out<=(others=>'Z');
		elsif(clk'event and clk='1') then
			data_out<=content(conv_integer(address));
		end if;
	end process;
end a_ROM_RGB;
