library ieee;
use ieee.std_logic_1164.all;

entity matrizRGB is port(
    clk: in std_logic;
    filas : out std_logic_vector(7 downto 0);
    rgb: out std_logic_vector(23 downto 0);
	f1,f2,f3,f4,f5,f6,f7,f8: in std_logic_vector(23 downto 0)
);
end matrizRGB;

architecture a_matrizRGB of matrizRGB is

signal temp_filas,temp_columna: std_logic_vector(7 downto 0):="00000001";
signal temp_rgb: std_logic_vector(23 downto 0):=(others=>'1');
signal c1,c2,c3,c4,c5,c6,c7,c8: std_logic_vector(23 downto 0):=(others=>'1');


begin

    process(clk)
    begin
        if(rising_edge(clk)) then
            case temp_filas is
                when "00000001"=>
                    temp_rgb <= c1;
                    temp_filas<="00000010";
                when "00000010"=>
                    temp_rgb <= c2;
                    temp_filas<="00000100";
                when "00000100"=>
                    temp_rgb <= c3;
                    temp_filas<="00001000";
                when "00001000"=>
                    temp_rgb <= c4;
                    temp_filas<="00010000";
                when "00010000"=>
                    temp_rgb <= c5;
                    temp_filas<="00100000";
                when "00100000"=>
                    temp_rgb <= c6;
                    temp_filas<="01000000";
                when "01000000"=>
                    temp_rgb <= c7;
                    temp_filas<="10000000";
                when "10000000"=>
                    temp_rgb <= c8;
                    temp_filas<="00000001";
                    
                    case temp_columna is
                        when "00000001"=>
                            c1<=f1(23)&f1(15)&f1(7)&"111111111111111111111";
                            c2<=f1(22)&f1(14)&f1(6)&"111111111111111111111";
                            c3<=f1(21)&f1(13)&f1(5)&"111111111111111111111";
                            c4<=f1(20)&f1(12)&f1(4)&"111111111111111111111";
                            c5<=f1(19)&f1(11)&f1(3)&"111111111111111111111";
                            c6<=f1(18)&f1(10)&f1(2)&"111111111111111111111";
                            c7<=f1(17)&f1(9)&f1(1)&"111111111111111111111";
                            c8<=f1(16)&f1(8)&f1(0)&"111111111111111111111";
                            temp_columna<="00000010";
                        when "00000010"=>
                            c1<="111"&f2(23)&f2(15)&f2(7)&"111111111111111111";
                            c2<="111"&f2(22)&f2(14)&f2(6)&"111111111111111111";
                            c3<="111"&f2(21)&f2(13)&f2(5)&"111111111111111111";
                            c4<="111"&f2(20)&f2(12)&f2(4)&"111111111111111111";
                            c5<="111"&f2(19)&f2(11)&f2(3)&"111111111111111111";
                            c6<="111"&f2(18)&f2(10)&f2(2)&"111111111111111111";
                            c7<="111"&f2(17)&f2(9)&f2(1)&"111111111111111111";
                            c8<="111"&f2(16)&f2(8)&f2(0)&"111111111111111111";
                            temp_columna<="00000100";
                        when "00000100"=>
                            c1<="111111"&f3(23)&f3(15)&f3(7)&"111111111111111";
                            c2<="111111"&f3(22)&f3(14)&f3(6)&"111111111111111";
                            c3<="111111"&f3(21)&f3(13)&f3(5)&"111111111111111";
                            c4<="111111"&f3(20)&f3(12)&f3(4)&"111111111111111";
                            c5<="111111"&f3(19)&f3(11)&f3(3)&"111111111111111";
                            c6<="111111"&f3(18)&f3(10)&f3(2)&"111111111111111";
                            c7<="111111"&f3(17)&f3(9)&f3(1)&"111111111111111";
                            c8<="111111"&f3(16)&f3(8)&f3(0)&"111111111111111";
                            temp_columna<="00001000";
                        when "00001000"=>
                            c1<="111111111"&f4(23)&f4(15)&f4(7)&"111111111111";
                            c2<="111111111"&f4(22)&f4(14)&f4(6)&"111111111111";
                            c3<="111111111"&f4(21)&f4(13)&f4(5)&"111111111111";
                            c4<="111111111"&f4(20)&f4(12)&f4(4)&"111111111111";
                            c5<="111111111"&f4(19)&f4(11)&f4(3)&"111111111111";
                            c6<="111111111"&f4(18)&f4(10)&f4(2)&"111111111111";
                            c7<="111111111"&f4(17)&f4(9)&f4(1)&"111111111111";
                            c8<="111111111"&f4(16)&f4(8)&f4(0)&"111111111111";
                            temp_columna<="00010000";
                        when "00010000"=>
                            c1<="111111111111"&f5(23)&f5(15)&f5(7)&"111111111";
                            c2<="111111111111"&f5(22)&f5(14)&f5(6)&"111111111";
                            c3<="111111111111"&f5(21)&f5(13)&f5(5)&"111111111";
                            c4<="111111111111"&f5(20)&f5(12)&f5(4)&"111111111";
                            c5<="111111111111"&f5(19)&f5(11)&f5(3)&"111111111";
                            c6<="111111111111"&f5(18)&f5(10)&f5(2)&"111111111";
                            c7<="111111111111"&f5(17)&f5(9)&f5(1)&"111111111";
                            c8<="111111111111"&f5(16)&f5(8)&f5(0)&"111111111";
                            temp_columna<="00100000";
                        when "00100000"=>
                            c1<="111111111111111"&f6(23)&f6(15)&f6(7)&"111111";
                            c2<="111111111111111"&f6(22)&f6(14)&f6(6)&"111111";
                            c3<="111111111111111"&f6(21)&f6(13)&f6(5)&"111111";
                            c4<="111111111111111"&f6(20)&f6(12)&f6(4)&"111111";
                            c5<="111111111111111"&f6(19)&f6(11)&f6(3)&"111111";
                            c6<="111111111111111"&f6(18)&f6(10)&f6(2)&"111111";
                            c7<="111111111111111"&f6(17)&f6(9)&f6(1)&"111111";
                            c8<="111111111111111"&f6(16)&f6(8)&f6(0)&"111111";
                            temp_columna<="01000000";
                        when "01000000"=>
                            c1<="111111111111111111"&f7(23)&f7(15)&f7(7)&"111";
                            c2<="111111111111111111"&f7(22)&f7(14)&f7(6)&"111";
                            c3<="111111111111111111"&f7(21)&f7(13)&f7(5)&"111";
                            c4<="111111111111111111"&f7(20)&f7(12)&f7(4)&"111";
                            c5<="111111111111111111"&f7(19)&f7(11)&f7(3)&"111";
                            c6<="111111111111111111"&f7(18)&f7(10)&f7(2)&"111";
                            c7<="111111111111111111"&f7(17)&f7(9)&f7(1)&"111";
                            c8<="111111111111111111"&f7(16)&f7(8)&f7(0)&"111";
                            temp_columna<="10000000";
                        when "10000000"=>
                            c1<="111111111111111111111"&f8(23)&f8(15)&f8(7);
                            c2<="111111111111111111111"&f8(22)&f8(14)&f8(6);
                            c3<="111111111111111111111"&f8(21)&f8(13)&f8(5);
                            c4<="111111111111111111111"&f8(20)&f8(12)&f8(4);
                            c5<="111111111111111111111"&f8(19)&f8(11)&f8(3);
                            c6<="111111111111111111111"&f8(18)&f8(10)&f8(2);
                            c7<="111111111111111111111"&f8(17)&f8(9)&f8(1);
                            c8<="111111111111111111111"&f8(16)&f8(8)&f8(0);
                            temp_columna<="00000001";
                        when others =>
                            temp_columna<="00000001";
                    end case;
                when others =>
                    temp_rgb <= (others => '1');
                    temp_filas<="00000001";
            end case;
        end if;
    end process;
    
    filas <= temp_filas;
    rgb<= temp_rgb;
    
end a_matrizRGB;
