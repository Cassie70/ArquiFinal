LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY bcdDisplay IS
	PORT(
	CLK,CLR: IN STD_LOGIC;
	E: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	DISPLAY:INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	
	);
END ENTITY bcdDisplay;

ARCHITECTURE behavior OF bcdDisplay IS
	CONSTANT DIG0: STD_LOGIC_VECTOR(6 DOWNTO 0):="0111111";
	CONSTANT DIG1: STD_LOGIC_VECTOR(6 DOWNTO 0):="0000110";
	CONSTANT DIG2: STD_LOGIC_VECTOR(6 DOWNTO 0):="1011011";
	CONSTANT DIG3: STD_LOGIC_VECTOR(6 DOWNTO 0):="1001111";
	CONSTANT DIG4: STD_LOGIC_VECTOR(6 DOWNTO 0):="1100110";
	CONSTANT DIG5: STD_LOGIC_VECTOR(6 DOWNTO 0):="1101101";
	CONSTANT DIG6: STD_LOGIC_VECTOR(6 DOWNTO 0):="1111101";
	CONSTANT DIG7: STD_LOGIC_VECTOR(6 DOWNTO 0):="0000111";
	CONSTANT DIG8: STD_LOGIC_VECTOR(6 DOWNTO 0):="1111111";
	CONSTANT DIG9: STD_LOGIC_VECTOR(6 DOWNTO 0):="1101111";
BEGIN
	PROCESS(CLK,CLR,DISPLAY,E)
BEGIN
	IF(CLR='1') THEN
	DISPLAY<=DIG0;
	ELSIF(CLK'EVENT AND CLK='1') THEN
		CASE E IS
			WHEN "0000"=>DISPLAY<=DIG0;
			WHEN "0001"=>DISPLAY<=DIG1;
			WHEN "0010"=>DISPLAY<=DIG2;
			WHEN "0011"=>DISPLAY<=DIG3;
			WHEN "0100"=>DISPLAY<=DIG4;
			WHEN "0101"=>DISPLAY<=DIG5;
			WHEN "0110"=>DISPLAY<=DIG6;
			WHEN "0111"=>DISPLAY<=DIG7;
			WHEN "1000"=>DISPLAY<=DIG8;
			WHEN OTHERS=>DISPLAY<=DIG9;
		END CASE;
	END IF;
	END PROCESS;
 END behavior;